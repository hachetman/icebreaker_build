// Convert 4bit numbers to 7 segments
module seven_seg_hex (
                      input [3:0] din,
                      output reg [6:0] dout
                      );
always @*
  case (din)
      4'h0: dout = 7'b 0111111;
      4'h1: dout = 7'b 0000110;
      4'h2: dout = 7'b 1011011;
      4'h3: dout = 7'b 1001111;
      4'h4: dout = 7'b 1100110;
      4'h5: dout = 7'b 1101101;
      4'h6: dout = 7'b 1111101;
      4'h7: dout = 7'b 0000111;
      4'h8: dout = 7'b 1111111;
      4'h9: dout = 7'b 1101111;
      4'hA: dout = 7'b 1110111;
      4'hB: dout = 7'b 1111100;
      4'hC: dout = 7'b 0111001;
      4'hD: dout = 7'b 1011110;
      4'hE: dout = 7'b 1111001;
      4'hF: dout = 7'b 1110001;
      default: dout = 7'b 1000000;
  endcase
endmodule
